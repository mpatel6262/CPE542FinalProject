`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 04/15/2024 02:47:29 PM
// Design Name: 
// Module Name: Matrix_Mult
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Matrix_Mult(

    );

    logic[127:0][31:0] memory;

    ProcessingElementMem PE1();

    PE_Controller PE1_cont();

endmodule
